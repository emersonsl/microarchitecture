
module processor (
	clk_clk,
	pio_0_external_connection_export,
	pio_1_external_connection_export);	

	input		clk_clk;
	output	[2:0]	pio_0_external_connection_export;
	input	[2:0]	pio_1_external_connection_export;
endmodule
